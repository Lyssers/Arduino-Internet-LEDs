PK   �:Y�<��*  ��    cirkitFile.json�}�n�ȑ�e�?���&����������mx�
,~��H���c�`h_�>�M������
2NJ�m`���yy2��<�ew����޷7���o�������0�������ߖ�����������w������Ǿ8��Mw��m�ա���U��r(t��E�iWH�����Z�/����N{���b{{1뿽����u}���ph��n��B��)%��l��e�D#�^�:/��y�y�s�y��w΃/9���Y�o~�o������?�\5����(����PL8&Ǒ%��5���{|1���;g+)*�W�]��C5��.���^��ԝa��]��`��p|Ǎ?�,>3�8d�qL	��o�����_�y��<nT%��ۦ1�����Z�uq\S8�D�*]�`5�y��<nUs�Ǎ`�d�0��I7��a2�	n2-,�J�$L��q�Pp����lS,��t�A����J�u�l=����Ӆ>��<ԍ.JQ[��9���ד�\Z2�E5�}�l��>v<5�9�JiI7���54�Zn<���B��s�X��㓉k£��(�&&*$�VH���9�tg����e��Ω҈�����L�l��4k�Ԗ�in��{���*�M:ǛI�AU)*!�o���*1t�1�(�\34�^�����y���O~�%S�Ji�2��5��nڦ�T%��9��:�7�)ɭY'�Lh�4�)I�&{Jj�7RymJV��gOIn���61�.�1躪V�EW��G�J��}�dUU�R��{Jr��$?Y�wJV�)I�&{J�&�J�hS�2�=%����,OG���g�XU1��f�xc<?	$�s|t�N`���������N`ѕ{������N`ѕ{������N`ѕ{������N`ѝ�A�Φ�[v�\�7��U�y���ezzo"�7��*��+��E�t=��Dxs<_�X��P�s��͉��i<�h9���E���?t]�.���� �V\[a�	0�q]�?p}��'���W`��k,,>�7�� �\ga�	0���7��zD��	0�q�ЪB��	0�q
���@��	0�q����^��	0�q�xi\`�	0�p�s)o�������o�,�/�����|���E��,>�7��\�`�	0�p�3|r�2Hp�������G��,>�7nI�\�`�	0�pCs�W��.����ك�\<Ip��'��[�[m��e��F���y����W��mD�u$�d~&l%�����ۃW6��]�|�!u-����9���k�3烘�0X�~�Gm{&���tk�3�![���-�m��_p^gm{&�$W(G
N�ܳ��fu�d��J�HÂϜ<�9yTz��x;�T�yD�3�n��q̽Q��yRs]�բB���s�[N��1O�
���s��(��d{��D-���RF��S�7���*�9M'����l#*�@w��\a���o4�f�ko+��(�T��ǋ*�J���SNymsP����y:�8زi�N�>8�����)����jн�����{�T׈a�J���x�wu_�J��1�v��;��B>uh�m��hu#]վy�l!��3����.�Nj�������w]��矮
���흰�4����{�����)��W5uQ[]){�Z-��.���|aܛҏP���S���(*cmQփ����pXwJ�t�CU�C��q�����hj����U��i�B����u��J�Tq~�6�w]Som�,�ޔ����{W��`����#>��\�H���`m#lg�N,�Nj��-{�v�oi^պ����Ӧ6�j��]�<�y�w�u�j�
a*�\W>R�,��۪���{'5_�64�!��w���LeuD��L�&D����w��S�Q%ӊQK�������T>OԾ�/��:u?~"������"a�۲��0p4^ģ!��M��oM�
��M��OK�|�<���?�C�p���0h6�C��E�Q<��Q��G�#s�5_x"��E�ȡx�h��"�P<z0��G5�G�!9��(QDz��g�(*=Z25,p�,E�1?ZBDJ�a�\�+3V
;㸅qܢ�p0?�,u�A�@��*����Q��}�;@b	z"�sG?5U����x���K�aq\*T̔
�I���a���[�s�pTd�	d�ϊ�$,��
�'X�S���F���B�K!&��h�g|i�X×�Dx T���u~|n�5� �[�u~�n��XC�P���-�V�~́5T�x`~n��XCuQ���+�V�~́5T�x`~�n����b<0?�	�
�k��j(��p�@���J�b<0?�	�
�k���'(��Q�D�?A9|��+ڈ$(�,ҷ�ʮ<uW ǉ7��m��+ڈ�(�,ҷyʯ,h#2�x�H��)����H���"}��˂6"O�7��m�R,ڈt)�,ҷyʱ,h#��x�H��)ɲ��H���"}��,˂6"��7�|���.˂6"��y�H�����.˂6���7��m�Wby�@�o��<uY��T�Y�o��eY�F�UA�6O]A�6��m��,�'9!O]�mDTo��<uY��UPL�S�EТ�"}��.DKAN�S��ЮWZXI��^��
���/�^�56}�+��޿�W?�Qb��z-T�����ʨ3���m�KE�Il�� ��0��p��EU��S�s6Ȭ"�`X�:��A{afbqxji��j�p�IT�MM,��lP8E<u1,VgYL�=����/]~zS�Hc:�EG,s���Ҡ�s��5>��B���u֫n�N9��ό�)_/�����eL`�.�e�o�^`r�/T��3~!
>�b|�
7.�*����:��V�r� +g�P�V�?�R� +g�P�V�b��8���Q�`�,��#��Y,T�G���X�� +g�P� V�b�JC���uD�Șz�z���5/�p�r�E`��'�R\�#� �r�E6Gz~��@��Q�?�O��w��}��?��6W��m:FA"���` ��Q0�d�(A2t� :
B�!�@����D CG�@"���@L��Em\؆�m�(K��L��-`�e�A0�	�,��,=b0�b��q���@&X��8��� ���˿q	8,�KXGYz�`��q	��(K��L�8.aqe�A0�	�%,��,�V��V#��h�0��@�U�_s`�B<�8B[�5ֈ` ��i#�U�_s`�B<�4B[�5ֈ` ��)#�U�_s`�B<�0B[�5ֈ` ���"�U�_s`�B<�,B[�5ֈ` ���"�U�_s`�b2�<W(�����\Y���f���Tv婻B	>�Y�o�^Y���f���S~eA��E�6O	�mL0n��<eX�1�@�Y�o�bY���f���S�eA��E�6OI�mL0n��<eY�1�@�Y䛅<uY�1�@�Y�o��eY���f����J,O]J���"}��.˂6&7��m��,ژ` �,ҷy�,hc��p�H��˲��	��"}��.˂6&7��m��,ژ` �,ҷy�2���|+����V��7�$�$o�[I��� ȷ��[�E0`���!�-�� 3�NGm��p8ulh�`  �aX�:O�E0`���A�-�� 3�N`l���XaX�β�,ȷ��rvB����V���,ȷr�/d�@���~!��U0�o�_���|+g�B�[9��` ��Y,d�@���q�*ȷrY0�o�,�` ��y�P�V�b!�bQ0�o�,�` ��Y,d�@����U0�o�|��
�`��}N��V��Y0p9JQ�V��]�`ࣕ_/��������������|y���?^5�������v������j��-Rt�_�Z��y��<�|�� �fv�S�gv�Xk�1���5����g��˶/*9Eߊ��md)Oo{��a�sbE��ܲ:g��q	�YK�x�1g�Wޘ3ëKuN\gau^�:g�y���HM�W���d�%�"�zONu�J�w��;��HC\���n����6���\4�/fVP4��A�H� f�^��A&wK� MZm�����ʕ�bh[Qh+DQپ�yn�z�;�)0�(����ά�&=����އ�=/.Nc�dE���'6�������-��j�C�����y��g�{�ٛ�dYy0Nߨ톺Х��ڛ-Z���uN��D�D�I��k*��%��ė:�^�Ay��Z�B�8o\ۺpM�M�eU@���Pzg{^$���ޓ��s�'�󝈝7ߓ�q�x���;k�%+_�̄q~Ȁ��Y]�A��TL,r���f���g�U�G�����[��|s�2�����r��#q��y���b�"� ]x��h��0y��Y�i^�;�E�B܆���#n�ʵ�@۰�k����*��0qkS��a���Ԧ�6>^��\�#n��=Փ/5���^{Q�1��|�8_Z���>�Ræ�r03��x�y�e"�L�� 4 �\�{���Ȝ�\�Ye��!���u_�d �f�A���}��O7�}s�����H�����F�	ëm\����|u����0����6Uծ��< ��<��7�s
�y�?����N-���Xu!�O���P�1��Q��"�E����X�v��?ρ��c%�����?d���?k��ᅎ��1�O��1 ��A Ρ,�x��(|�S)|��)|�3*����
��
��
�>�_ɵ���/��7s�|	0����0 �g�0 �G�����p���q�����Gi�a=q�0?Fѿ��b�7�m�����ԍ�®� ���q���B*n�=�#�X�e� �W=dHH�^��!�"�$"�@"�\"�x" �r�ƹc� ��3ϒ�:4�8;�8B
�D��\;;^5N�#�k�j@Bn@B�q�;Y���g�$؅K��4���}N�(�C�R�_�!�|�>a��yj�5OEg�܊�[QC@p+j��܆70���o`�Ҋ�������!��w�_��&�G{���o�Q)H@F�^����dQ�F)5WG�L��")��]#W�D ��ĸ�l��Yd��/g �3o�Gok(��Ɔ�+�XO�9G����>�*ݓ�E=Q�'�z��O�=�T=��{*��>���K��,��|!��E/���a��6��[Y6ɥ��ıMz�,�uGr[�+���p�n�Z�G�#�N�ל� �&�G��M|���1ya���bN|M'��_�	�/���{�8v�ɧ����}s�����a8v������v��9���<�omZD,��Y+B����%3䏟���@�3�W��XsUD,����N��bɌPN��b�_�O@�b>����Œp+8C�%�I]�	Z,�e@�g����yz091�ML����1U>��1)�g"nF�d/����
nQ(�0Ϟ�I����yl�q>��i�>j5���L%�~�L��XLa��$�J Dy����9���u��d�+��3��$��P�{��dbۘVm�)�nfἅnq4Ʌ�q�*���	,�*Q ���r�1�w�"D���2�+��N��	0>��'��?,>�W��
�?,>�W�5��?,>�W���?,>�w"B	�]~��-�W�p�����tg��J���2o���:�,2ى�+B��ۯ��ϸ��W\��.7W��1�7�|#ߡ�}�`�%���"F��0B�F8��B�]ɀ
4���ڇ�j�P��o��>DW4`��p|��!�Lh��p|I��!�6h��p|���!� h��p|9��!�
h��0<�
5�Y�F�)`��Y��	|UB��ea�;5��!���l��E��0B�Fj%@b|�.[�CY���6<����0�q���*�P����>DW1`��0��Z��ĳ�q)��#?O5��!��9�p��S��we�`��Z�)f�`G��.o�[����ms+�;?W��h�l�\�>����]lzr���Yk��P�^k �Ǽ� ������D�Q��S\&�G��21���� ���M��c/r�)!}E���id?{J��f�K[ť�Z�m��C[U�pC��/M�(o�l��e�D#�J�!'�����(�"����$s���	�@g+)*�W�]��C5����1��� ugb�Kd$s�%r����2�$s�%�t�4���0Z�B��.�k
'����P�k"��� ���&N��d.⻄p �\�w�8�ke�5Em�.���<ԍ.|�i���P�6��Ȓ�E|�Y���w"1gI�Ν|~2���H�`��և U��E���5Z�T�TP��/�ۃ-���t1�����n��JkJ��;��?��B���1��C����ή�Z��3f��'�_z�Za۾+Z��BW�o�*[�f�L��������/�oz|T���_��'��
���흰�4K���/���C��зR�;�j��*�R���Z֝]�����7��Je�*�:QT�ڢ�W����8����U���Ʃڷ�ˢ�}�b:3T}?��UK���/��k?CmW�����m￦2���gNY�)��'�_�_�y�\]�>s����Ԫ�6�v���R�����e�ڮ�M���Z�މ�ԦS�����'�_��i]�کB�ʷ�U_4'��<�ꤲz��I��M�vY`�B����ժ������|D}���ۮ����b���|�z������j��H)������e7��y�w���۽��=6�H��y#��1o},F�<s�=��S�=�OSJ6�yS�8-�NK�S�>��4� O�x=͕�C�o'��I�z��Vc_�~�%�c!|ߐR�DR�xCBmH�����%#;i@I�NPr���$��Y�IJpҀ��>i@yО4�<OPe�Gx:���7�D٠%Z��0������18��c���66���^rVvB<%o���s�= �7ɼ7�*Z��N�^��܋���L�$rB�JY��$�C\�c��D�X�8�̹�����5S��E�T	<ĥC�*����ar��n�f��2�X�!�g3�("�Q� �b,P$4�ԣ�����#����b<���9>�D�<o� � D�����{h�ԣ���.>����oam����iwSs��V��Qpw���K�m��`��-�^���&g�5�^݊�R$g�6�;Ž;�9k�������� �A�j��o���r�p������xSp;�@}��!�&����-2&8_�d�F�|��������9�W�����������3ơ�O��Oe��|�I�?���T��~�I�?���L��}�Ɇ?���\�S��S�T?�T?��[�=�Ϟ
]%�!B��G���#��#"t�xt�}"}"B��G���+��+"t�xt��"�"C���\�]>�L�>��~��_�_d����E>����󿹺�?�;��������~KUW��I?��`�?�Cq(USXW��7��5ro�^��|����R��~��M��OAU>��|w��+]�?}��ȥ���y�������2�շ�7����~z������_c��.���������u�������5W�����o������Ɩ�Z��G�}����w�Ow?����������]���o�rywy��?��m�ߟ.o�n���߀����OC����o��<���?����~���
@���L�����;僪̻J*Q��9Z;!܅(�wu�5B?N»y�{oa��k�r8��[��uea�?m�u�`��g����}s�ې^W_�nn/�86G`;?�~t/o۫�ad?(+ߙQ��/>(��\?��.�����_/��t�����K{w�,މw��A_���)~�<5�;?���=�U.7H;����<�}���|)n���k� %���UF8
�Ä����.������䐪;]��SN�mє�PT��������M�@�BI��9�Z_�z�D��L�"�TY%��d�l��md�������5a�mt��J�I�V��J]hq���u��-į3�v�"ړD{%͞�i��#ڳD{�h/dQ��2��u�ů��.�e������B�Ư^�5��>5|���M"H�	�	#�������y��{�$���ϸa&e��e*�V<q��'nX���-���.�ȟLw�i���yv�Ӱ�is��p�������臨�������E]�NԵ��}nV�b\b���U;��!w7?_?!z��	���ѧGw�M��I3�U�N�5���g9�����?�%}�K����O���7~�Ms��-�_��Ҝ����?��B5�O#J����BzR��Yغ�jSJ��Nz�c�CӨ�Խ�	mc�^�Ak�V�i�,&�&�XT�)zY_(]��O����r�����l�~e���Ӆ"i/��a�TU�]��沜��˅�j��_���F�(�.T]��.�3e)�֊�c�ɒ-��Ϲ:J��_��%Y�>��X�r�K:�-Ϙ��B���W�~I�B��gȤ�v�b�.s��2�Kb�~W	�5�]�]�c��זּ�U�w��Kc�	Ѝ46)��4��hl�=笐�~;��N�)�7&.�H�釯<��xl|�-M�	��z����b�i��,�+������Y:l������$�-��`��:��+ǿl�k0�I�#9b9�����8~al�фGj�6ζ$�5��˾���"�l�����'�9m�x�5���-�m���Zc�=v&|/�]m�S'{ZD�Z�3.TVE_�X#ۢ�A����৫�=+ʦ��QgմSz�+���g�����*Q*y|�pl��ָ��譇-y֠�E���v�w�����~���?���|��;��t��3$�2��(g�F=P��oƍ��OT�0a�q<?t��1��|������x�k:��~W�0s���|���8��i����~ܭ6E��]i�41�>o���ֽ�ۦ����|~���������/*����w~̮nn�۽�n�[?u�a�nw�����������w�Oɶ�^�E��Up�L�6?��,���ӡ�OF�d���~��������q���w�}����a�v��O�nŻ�o��)��H�?ݫ4^p1�c:��*Q��U�����WϚ9�o���Q@䣀S@ (PEw:7���7K��aNJ�eJ@�����>�!�i=�(N�ap8A.F����1�DĈz>����n��#�8�2�A�z�Ut
�%<Y�$
�$V�Q@�)�*�������j�U�La�S��(�1
0Q@��������U�E��@�z��)����8�f�Uo�\=蜔���z!1��J��E�F�a�� #2�#�B8l�ٯ�n�*z�P
�,V$
�$��Q��S`T&\tz�-WQ) �%c��@�d�S �,�v��Âtիf
�������q�`��Xy$����p��%��YIO#�y	cb�����J*a45�"��E�G72Rb���
��8!���_��닂�������$X�aV&	ttx��p՚F�^a�Uf��e2�`�2�
�L�h����^��m���A��$X�м+�.>�Ն��.	�_V�J
x���L����_�/��(h/#h���H�o#V`eƉ:�n�U�8��M�/�`�Ġ1��{b��	*0*DЮ�Ĥ&�lm|���Q�Մ��f�������0k?8���&�y���q2�MS�3{ky��H<QHQ�c����3~x���!~�/�sg���T;��Yv%Y�I$ػ��������p���#훊Yy �<X�u-N�N&���(�*��nB���Õ�G��;�YQ����h�i�\�V��G�76lZ�����>��Zq1T��\�&mŊ��׌,0蔠BL�������/���Iڧ{��V`eF���~>�V\V$�u��j*4	h�3��K����l�(������Q��k����< G�Xy� 1���Ԛ��k�E����3�Bg("���C�Ԍ�pQ�`y+$Y�������*">�O
�~5o�C�N9�_(R�"E<3���1���B���霑���H��S1"�UĜb4����Lrl�7�#L0	6���� ��9��ޥ��ْg���Ϣ϶JBR�:�v:�^de�ݤ���]��[*L7�5��.R�Ȼ�2#X|s������P�����t�s3�0�e$��|�8����� ]�b�:s�gi{�Vf����MB/���R�:w�8�MK��c!����&'��̘�J~��Hu�w����7�Y�w���f���D2OH�?�S����r����zM�-m��L�,;�%�E^H�ߋ1���9Kp�RgiU~+�0��)!ĉ/�ωC�*N�y�B���8K��[i��8g��9��$����%hW%�5'qˀi[�zt�K;Mz��3�U�����x�3à���2���7�%O�����Iw�g���L��V�5[�U�I��C�隅_gO����YgPN�C�(��y�\���Yڸ���Yxsv3���$�)�҆tQ�[�|�x�6�J���]3�Fڨ;OtZOA�(��9m�����\^]�a��澿�l��v�G&�M�q�?}������ꛛ�~��t7�����~��PK
   �:Y�<��*  ��                  cirkitFile.jsonPK      =   ?*    